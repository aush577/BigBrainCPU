module ewb_datapath
(
  input clk,
  input rst
);


endmodule : ewb_datapath
