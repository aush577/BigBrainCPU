module btb();

//branch target buffer




endmodule