module ewb_control
(
  input clk,
  input rst
);


endmodule : ewb_control
