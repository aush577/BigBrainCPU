module datapath (

);


endmodule : datapth
